
module system (
	clk_clk,
	reset_reset_n,
	ws2812_controller_0_conduit_end_regout);	

	input		clk_clk;
	input		reset_reset_n;
	output		ws2812_controller_0_conduit_end_regout;
endmodule
