
module N_leds (
	clk_clk,
	reset_reset_n,
	n_leds_controller_0_conduit_end_regout);	

	input		clk_clk;
	input		reset_reset_n;
	output		n_leds_controller_0_conduit_end_regout;
endmodule
